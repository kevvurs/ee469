this file is to test the git push shit