module fowarding (
);